/// Математические функции и константы
package math;

/// Математические функции и константы
class math;

    /// Число π
    static const real pi = 3.1415926535897931;

    /// Число е (число Эйлера)
    static const real e = 2.7182818284590451;

endclass

endpackage