// Таблица SIN (10'b -> 16'b)
/*
    SVERDLOVSK
    system verilog library

    Neveroff M.V.
    2025
*/

module ram_sin (
    i_val,
    o_val
    );

    input  [15:0] i_val;
    output [15:0] o_val;

    always_comb begin
        o_val = 'h0000;

        case (i_val[15:6])
            'h000: o_val = 'h7FFF;
            'h001: o_val = 'h80C8;
            'h002: o_val = 'h8191;
            'h003: o_val = 'h825A;
            'h004: o_val = 'h8323;
            'h005: o_val = 'h83EC;
            'h006: o_val = 'h84B5;
            'h007: o_val = 'h857E;
            'h008: o_val = 'h8647;
            'h009: o_val = 'h8710;
            'h00A: o_val = 'h87D8;
            'h00B: o_val = 'h88A1;
            'h00C: o_val = 'h896A;
            'h00D: o_val = 'h8A32;
            'h00E: o_val = 'h8AFA;
            'h00F: o_val = 'h8BC3;
            'h010: o_val = 'h8C8B;
            'h011: o_val = 'h8D53;
            'h012: o_val = 'h8E1B;
            'h013: o_val = 'h8EE2;
            'h014: o_val = 'h8FAA;
            'h015: o_val = 'h9072;
            'h016: o_val = 'h9139;
            'h017: o_val = 'h9200;
            'h018: o_val = 'h92C7;
            'h019: o_val = 'h938E;
            'h01A: o_val = 'h9454;
            'h01B: o_val = 'h951B;
            'h01C: o_val = 'h95E1;
            'h01D: o_val = 'h96A7;
            'h01E: o_val = 'h976D;
            'h01F: o_val = 'h9832;
            'h020: o_val = 'h98F8;
            'h021: o_val = 'h99BD;
            'h022: o_val = 'h9A82;
            'h023: o_val = 'h9B46;
            'h024: o_val = 'h9C0A;
            'h025: o_val = 'h9CCE;
            'h026: o_val = 'h9D92;
            'h027: o_val = 'h9E56;
            'h028: o_val = 'h9F19;
            'h029: o_val = 'h9FDC;
            'h02A: o_val = 'hA09E;
            'h02B: o_val = 'hA161;
            'h02C: o_val = 'hA223;
            'h02D: o_val = 'hA2E4;
            'h02E: o_val = 'hA3A5;
            'h02F: o_val = 'hA466;
            'h030: o_val = 'hA527;
            'h031: o_val = 'hA5E7;
            'h032: o_val = 'hA6A7;
            'h033: o_val = 'hA766;
            'h034: o_val = 'hA826;
            'h035: o_val = 'hA8E4;
            'h036: o_val = 'hA9A3;
            'h037: o_val = 'hAA61;
            'h038: o_val = 'hAB1E;
            'h039: o_val = 'hABDB;
            'h03A: o_val = 'hAC98;
            'h03B: o_val = 'hAD54;
            'h03C: o_val = 'hAE10;
            'h03D: o_val = 'hAECB;
            'h03E: o_val = 'hAF86;
            'h03F: o_val = 'hB041;
            'h040: o_val = 'hB0FB;
            'h041: o_val = 'hB1B4;
            'h042: o_val = 'hB26D;
            'h043: o_val = 'hB326;
            'h044: o_val = 'hB3DE;
            'h045: o_val = 'hB495;
            'h046: o_val = 'hB54C;
            'h047: o_val = 'hB603;
            'h048: o_val = 'hB6B9;
            'h049: o_val = 'hB76E;
            'h04A: o_val = 'hB823;
            'h04B: o_val = 'hB8D8;
            'h04C: o_val = 'hB98C;
            'h04D: o_val = 'hBA3F;
            'h04E: o_val = 'hBAF2;
            'h04F: o_val = 'hBBA4;
            'h050: o_val = 'hBC55;
            'h051: o_val = 'hBD07;
            'h052: o_val = 'hBDB7;
            'h053: o_val = 'hBE67;
            'h054: o_val = 'hBF16;
            'h055: o_val = 'hBFC5;
            'h056: o_val = 'hC073;
            'h057: o_val = 'hC120;
            'h058: o_val = 'hC1CD;
            'h059: o_val = 'hC279;
            'h05A: o_val = 'hC324;
            'h05B: o_val = 'hC3CF;
            'h05C: o_val = 'hC47A;
            'h05D: o_val = 'hC523;
            'h05E: o_val = 'hC5CC;
            'h05F: o_val = 'hC674;
            'h060: o_val = 'hC71C;
            'h061: o_val = 'hC7C2;
            'h062: o_val = 'hC869;
            'h063: o_val = 'hC90E;
            'h064: o_val = 'hC9B3;
            'h065: o_val = 'hCA57;
            'h066: o_val = 'hCAFA;
            'h067: o_val = 'hCB9D;
            'h068: o_val = 'hCC3F;
            'h069: o_val = 'hCCE0;
            'h06A: o_val = 'hCD80;
            'h06B: o_val = 'hCE20;
            'h06C: o_val = 'hCEBF;
            'h06D: o_val = 'hCF5D;
            'h06E: o_val = 'hCFFA;
            'h06F: o_val = 'hD097;
            'h070: o_val = 'hD132;
            'h071: o_val = 'hD1CE;
            'h072: o_val = 'hD268;
            'h073: o_val = 'hD301;
            'h074: o_val = 'hD39A;
            'h075: o_val = 'hD432;
            'h076: o_val = 'hD4C9;
            'h077: o_val = 'hD55F;
            'h078: o_val = 'hD5F4;
            'h079: o_val = 'hD689;
            'h07A: o_val = 'hD71D;
            'h07B: o_val = 'hD7AF;
            'h07C: o_val = 'hD842;
            'h07D: o_val = 'hD8D3;
            'h07E: o_val = 'hD963;
            'h07F: o_val = 'hD9F3;
            'h080: o_val = 'hDA81;
            'h081: o_val = 'hDB0F;
            'h082: o_val = 'hDB9C;
            'h083: o_val = 'hDC28;
            'h084: o_val = 'hDCB3;
            'h085: o_val = 'hDD3D;
            'h086: o_val = 'hDDC6;
            'h087: o_val = 'hDE4F;
            'h088: o_val = 'hDED6;
            'h089: o_val = 'hDF5D;
            'h08A: o_val = 'hDFE2;
            'h08B: o_val = 'hE067;
            'h08C: o_val = 'hE0EB;
            'h08D: o_val = 'hE16E;
            'h08E: o_val = 'hE1F0;
            'h08F: o_val = 'hE271;
            'h090: o_val = 'hE2F1;
            'h091: o_val = 'hE370;
            'h092: o_val = 'hE3EE;
            'h093: o_val = 'hE46B;
            'h094: o_val = 'hE4E7;
            'h095: o_val = 'hE562;
            'h096: o_val = 'hE5DD;
            'h097: o_val = 'hE656;
            'h098: o_val = 'hE6CE;
            'h099: o_val = 'hE745;
            'h09A: o_val = 'hE7BC;
            'h09B: o_val = 'hE831;
            'h09C: o_val = 'hE8A5;
            'h09D: o_val = 'hE918;
            'h09E: o_val = 'hE98B;
            'h09F: o_val = 'hE9FC;
            'h0A0: o_val = 'hEA6C;
            'h0A1: o_val = 'hEADB;
            'h0A2: o_val = 'hEB4A;
            'h0A3: o_val = 'hEBB7;
            'h0A4: o_val = 'hEC23;
            'h0A5: o_val = 'hEC8E;
            'h0A6: o_val = 'hECF8;
            'h0A7: o_val = 'hED61;
            'h0A8: o_val = 'hEDC9;
            'h0A9: o_val = 'hEE2F;
            'h0AA: o_val = 'hEE95;
            'h0AB: o_val = 'hEEFA;
            'h0AC: o_val = 'hEF5E;
            'h0AD: o_val = 'hEFC0;
            'h0AE: o_val = 'hF022;
            'h0AF: o_val = 'hF082;
            'h0B0: o_val = 'hF0E1;
            'h0B1: o_val = 'hF140;
            'h0B2: o_val = 'hF19D;
            'h0B3: o_val = 'hF1F9;
            'h0B4: o_val = 'hF254;
            'h0B5: o_val = 'hF2AE;
            'h0B6: o_val = 'hF306;
            'h0B7: o_val = 'hF35E;
            'h0B8: o_val = 'hF3B4;
            'h0B9: o_val = 'hF40A;
            'h0BA: o_val = 'hF45E;
            'h0BB: o_val = 'hF4B1;
            'h0BC: o_val = 'hF503;
            'h0BD: o_val = 'hF554;
            'h0BE: o_val = 'hF5A4;
            'h0BF: o_val = 'hF5F3;
            'h0C0: o_val = 'hF640;
            'h0C1: o_val = 'hF68D;
            'h0C2: o_val = 'hF6D8;
            'h0C3: o_val = 'hF722;
            'h0C4: o_val = 'hF76B;
            'h0C5: o_val = 'hF7B3;
            'h0C6: o_val = 'hF7F9;
            'h0C7: o_val = 'hF83F;
            'h0C8: o_val = 'hF883;
            'h0C9: o_val = 'hF8C6;
            'h0CA: o_val = 'hF908;
            'h0CB: o_val = 'hF949;
            'h0CC: o_val = 'hF989;
            'h0CD: o_val = 'hF9C7;
            'h0CE: o_val = 'hFA04;
            'h0CF: o_val = 'hFA41;
            'h0D0: o_val = 'hFA7C;
            'h0D1: o_val = 'hFAB5;
            'h0D2: o_val = 'hFAEE;
            'h0D3: o_val = 'hFB25;
            'h0D4: o_val = 'hFB5C;
            'h0D5: o_val = 'hFB91;
            'h0D6: o_val = 'hFBC4;
            'h0D7: o_val = 'hFBF7;
            'h0D8: o_val = 'hFC28;
            'h0D9: o_val = 'hFC59;
            'h0DA: o_val = 'hFC88;
            'h0DB: o_val = 'hFCB6;
            'h0DC: o_val = 'hFCE2;
            'h0DD: o_val = 'hFD0E;
            'h0DE: o_val = 'hFD38;
            'h0DF: o_val = 'hFD61;
            'h0E0: o_val = 'hFD89;
            'h0E1: o_val = 'hFDB0;
            'h0E2: o_val = 'hFDD5;
            'h0E3: o_val = 'hFDF9;
            'h0E4: o_val = 'hFE1C;
            'h0E5: o_val = 'hFE3E;
            'h0E6: o_val = 'hFE5E;
            'h0E7: o_val = 'hFE7E;
            'h0E8: o_val = 'hFE9C;
            'h0E9: o_val = 'hFEB9;
            'h0EA: o_val = 'hFED4;
            'h0EB: o_val = 'hFEEF;
            'h0EC: o_val = 'hFF08;
            'h0ED: o_val = 'hFF20;
            'h0EE: o_val = 'hFF37;
            'h0EF: o_val = 'hFF4C;
            'h0F0: o_val = 'hFF61;
            'h0F1: o_val = 'hFF74;
            'h0F2: o_val = 'hFF86;
            'h0F3: o_val = 'hFF96;
            'h0F4: o_val = 'hFFA6;
            'h0F5: o_val = 'hFFB4;
            'h0F6: o_val = 'hFFC1;
            'h0F7: o_val = 'hFFCD;
            'h0F8: o_val = 'hFFD7;
            'h0F9: o_val = 'hFFE0;
            'h0FA: o_val = 'hFFE8;
            'h0FB: o_val = 'hFFEF;
            'h0FC: o_val = 'hFFF5;
            'h0FD: o_val = 'hFFF9;
            'h0FE: o_val = 'hFFFC;
            'h0FF: o_val = 'hFFFE;
            'h100: o_val = 'hFFFF;
            'h101: o_val = 'hFFFE;
            'h102: o_val = 'hFFFC;
            'h103: o_val = 'hFFF9;
            'h104: o_val = 'hFFF5;
            'h105: o_val = 'hFFEF;
            'h106: o_val = 'hFFE8;
            'h107: o_val = 'hFFE0;
            'h108: o_val = 'hFFD7;
            'h109: o_val = 'hFFCD;
            'h10A: o_val = 'hFFC1;
            'h10B: o_val = 'hFFB4;
            'h10C: o_val = 'hFFA6;
            'h10D: o_val = 'hFF96;
            'h10E: o_val = 'hFF86;
            'h10F: o_val = 'hFF74;
            'h110: o_val = 'hFF61;
            'h111: o_val = 'hFF4C;
            'h112: o_val = 'hFF37;
            'h113: o_val = 'hFF20;
            'h114: o_val = 'hFF08;
            'h115: o_val = 'hFEEF;
            'h116: o_val = 'hFED4;
            'h117: o_val = 'hFEB9;
            'h118: o_val = 'hFE9C;
            'h119: o_val = 'hFE7E;
            'h11A: o_val = 'hFE5E;
            'h11B: o_val = 'hFE3E;
            'h11C: o_val = 'hFE1C;
            'h11D: o_val = 'hFDF9;
            'h11E: o_val = 'hFDD5;
            'h11F: o_val = 'hFDB0;
            'h120: o_val = 'hFD89;
            'h121: o_val = 'hFD61;
            'h122: o_val = 'hFD38;
            'h123: o_val = 'hFD0E;
            'h124: o_val = 'hFCE2;
            'h125: o_val = 'hFCB6;
            'h126: o_val = 'hFC88;
            'h127: o_val = 'hFC59;
            'h128: o_val = 'hFC28;
            'h129: o_val = 'hFBF7;
            'h12A: o_val = 'hFBC4;
            'h12B: o_val = 'hFB91;
            'h12C: o_val = 'hFB5C;
            'h12D: o_val = 'hFB25;
            'h12E: o_val = 'hFAEE;
            'h12F: o_val = 'hFAB5;
            'h130: o_val = 'hFA7C;
            'h131: o_val = 'hFA41;
            'h132: o_val = 'hFA04;
            'h133: o_val = 'hF9C7;
            'h134: o_val = 'hF989;
            'h135: o_val = 'hF949;
            'h136: o_val = 'hF908;
            'h137: o_val = 'hF8C6;
            'h138: o_val = 'hF883;
            'h139: o_val = 'hF83F;
            'h13A: o_val = 'hF7F9;
            'h13B: o_val = 'hF7B3;
            'h13C: o_val = 'hF76B;
            'h13D: o_val = 'hF722;
            'h13E: o_val = 'hF6D8;
            'h13F: o_val = 'hF68D;
            'h140: o_val = 'hF640;
            'h141: o_val = 'hF5F3;
            'h142: o_val = 'hF5A4;
            'h143: o_val = 'hF554;
            'h144: o_val = 'hF503;
            'h145: o_val = 'hF4B1;
            'h146: o_val = 'hF45E;
            'h147: o_val = 'hF40A;
            'h148: o_val = 'hF3B4;
            'h149: o_val = 'hF35E;
            'h14A: o_val = 'hF306;
            'h14B: o_val = 'hF2AE;
            'h14C: o_val = 'hF254;
            'h14D: o_val = 'hF1F9;
            'h14E: o_val = 'hF19D;
            'h14F: o_val = 'hF140;
            'h150: o_val = 'hF0E1;
            'h151: o_val = 'hF082;
            'h152: o_val = 'hF022;
            'h153: o_val = 'hEFC0;
            'h154: o_val = 'hEF5E;
            'h155: o_val = 'hEEFA;
            'h156: o_val = 'hEE95;
            'h157: o_val = 'hEE2F;
            'h158: o_val = 'hEDC9;
            'h159: o_val = 'hED61;
            'h15A: o_val = 'hECF8;
            'h15B: o_val = 'hEC8E;
            'h15C: o_val = 'hEC23;
            'h15D: o_val = 'hEBB7;
            'h15E: o_val = 'hEB4A;
            'h15F: o_val = 'hEADB;
            'h160: o_val = 'hEA6C;
            'h161: o_val = 'hE9FC;
            'h162: o_val = 'hE98B;
            'h163: o_val = 'hE918;
            'h164: o_val = 'hE8A5;
            'h165: o_val = 'hE831;
            'h166: o_val = 'hE7BC;
            'h167: o_val = 'hE745;
            'h168: o_val = 'hE6CE;
            'h169: o_val = 'hE656;
            'h16A: o_val = 'hE5DD;
            'h16B: o_val = 'hE562;
            'h16C: o_val = 'hE4E7;
            'h16D: o_val = 'hE46B;
            'h16E: o_val = 'hE3EE;
            'h16F: o_val = 'hE370;
            'h170: o_val = 'hE2F1;
            'h171: o_val = 'hE271;
            'h172: o_val = 'hE1F0;
            'h173: o_val = 'hE16E;
            'h174: o_val = 'hE0EB;
            'h175: o_val = 'hE067;
            'h176: o_val = 'hDFE2;
            'h177: o_val = 'hDF5D;
            'h178: o_val = 'hDED6;
            'h179: o_val = 'hDE4F;
            'h17A: o_val = 'hDDC6;
            'h17B: o_val = 'hDD3D;
            'h17C: o_val = 'hDCB3;
            'h17D: o_val = 'hDC28;
            'h17E: o_val = 'hDB9C;
            'h17F: o_val = 'hDB0F;
            'h180: o_val = 'hDA81;
            'h181: o_val = 'hD9F3;
            'h182: o_val = 'hD963;
            'h183: o_val = 'hD8D3;
            'h184: o_val = 'hD842;
            'h185: o_val = 'hD7AF;
            'h186: o_val = 'hD71D;
            'h187: o_val = 'hD689;
            'h188: o_val = 'hD5F4;
            'h189: o_val = 'hD55F;
            'h18A: o_val = 'hD4C9;
            'h18B: o_val = 'hD432;
            'h18C: o_val = 'hD39A;
            'h18D: o_val = 'hD301;
            'h18E: o_val = 'hD268;
            'h18F: o_val = 'hD1CE;
            'h190: o_val = 'hD132;
            'h191: o_val = 'hD097;
            'h192: o_val = 'hCFFA;
            'h193: o_val = 'hCF5D;
            'h194: o_val = 'hCEBF;
            'h195: o_val = 'hCE20;
            'h196: o_val = 'hCD80;
            'h197: o_val = 'hCCE0;
            'h198: o_val = 'hCC3F;
            'h199: o_val = 'hCB9D;
            'h19A: o_val = 'hCAFA;
            'h19B: o_val = 'hCA57;
            'h19C: o_val = 'hC9B3;
            'h19D: o_val = 'hC90E;
            'h19E: o_val = 'hC869;
            'h19F: o_val = 'hC7C2;
            'h1A0: o_val = 'hC71C;
            'h1A1: o_val = 'hC674;
            'h1A2: o_val = 'hC5CC;
            'h1A3: o_val = 'hC523;
            'h1A4: o_val = 'hC47A;
            'h1A5: o_val = 'hC3CF;
            'h1A6: o_val = 'hC324;
            'h1A7: o_val = 'hC279;
            'h1A8: o_val = 'hC1CD;
            'h1A9: o_val = 'hC120;
            'h1AA: o_val = 'hC073;
            'h1AB: o_val = 'hBFC5;
            'h1AC: o_val = 'hBF16;
            'h1AD: o_val = 'hBE67;
            'h1AE: o_val = 'hBDB7;
            'h1AF: o_val = 'hBD07;
            'h1B0: o_val = 'hBC55;
            'h1B1: o_val = 'hBBA4;
            'h1B2: o_val = 'hBAF2;
            'h1B3: o_val = 'hBA3F;
            'h1B4: o_val = 'hB98C;
            'h1B5: o_val = 'hB8D8;
            'h1B6: o_val = 'hB823;
            'h1B7: o_val = 'hB76E;
            'h1B8: o_val = 'hB6B9;
            'h1B9: o_val = 'hB603;
            'h1BA: o_val = 'hB54C;
            'h1BB: o_val = 'hB495;
            'h1BC: o_val = 'hB3DE;
            'h1BD: o_val = 'hB326;
            'h1BE: o_val = 'hB26D;
            'h1BF: o_val = 'hB1B4;
            'h1C0: o_val = 'hB0FB;
            'h1C1: o_val = 'hB041;
            'h1C2: o_val = 'hAF86;
            'h1C3: o_val = 'hAECB;
            'h1C4: o_val = 'hAE10;
            'h1C5: o_val = 'hAD54;
            'h1C6: o_val = 'hAC98;
            'h1C7: o_val = 'hABDB;
            'h1C8: o_val = 'hAB1E;
            'h1C9: o_val = 'hAA61;
            'h1CA: o_val = 'hA9A3;
            'h1CB: o_val = 'hA8E4;
            'h1CC: o_val = 'hA826;
            'h1CD: o_val = 'hA766;
            'h1CE: o_val = 'hA6A7;
            'h1CF: o_val = 'hA5E7;
            'h1D0: o_val = 'hA527;
            'h1D1: o_val = 'hA466;
            'h1D2: o_val = 'hA3A5;
            'h1D3: o_val = 'hA2E4;
            'h1D4: o_val = 'hA223;
            'h1D5: o_val = 'hA161;
            'h1D6: o_val = 'hA09E;
            'h1D7: o_val = 'h9FDC;
            'h1D8: o_val = 'h9F19;
            'h1D9: o_val = 'h9E56;
            'h1DA: o_val = 'h9D92;
            'h1DB: o_val = 'h9CCE;
            'h1DC: o_val = 'h9C0A;
            'h1DD: o_val = 'h9B46;
            'h1DE: o_val = 'h9A82;
            'h1DF: o_val = 'h99BD;
            'h1E0: o_val = 'h98F8;
            'h1E1: o_val = 'h9832;
            'h1E2: o_val = 'h976D;
            'h1E3: o_val = 'h96A7;
            'h1E4: o_val = 'h95E1;
            'h1E5: o_val = 'h951B;
            'h1E6: o_val = 'h9454;
            'h1E7: o_val = 'h938E;
            'h1E8: o_val = 'h92C7;
            'h1E9: o_val = 'h9200;
            'h1EA: o_val = 'h9139;
            'h1EB: o_val = 'h9072;
            'h1EC: o_val = 'h8FAA;
            'h1ED: o_val = 'h8EE2;
            'h1EE: o_val = 'h8E1B;
            'h1EF: o_val = 'h8D53;
            'h1F0: o_val = 'h8C8B;
            'h1F1: o_val = 'h8BC3;
            'h1F2: o_val = 'h8AFA;
            'h1F3: o_val = 'h8A32;
            'h1F4: o_val = 'h896A;
            'h1F5: o_val = 'h88A1;
            'h1F6: o_val = 'h87D8;
            'h1F7: o_val = 'h8710;
            'h1F8: o_val = 'h8647;
            'h1F9: o_val = 'h857E;
            'h1FA: o_val = 'h84B5;
            'h1FB: o_val = 'h83EC;
            'h1FC: o_val = 'h8323;
            'h1FD: o_val = 'h825A;
            'h1FE: o_val = 'h8191;
            'h1FF: o_val = 'h80C8;
            'h200: o_val = 'h7FFF;
            'h201: o_val = 'h7F36;
            'h202: o_val = 'h7E6D;
            'h203: o_val = 'h7DA4;
            'h204: o_val = 'h7CDB;
            'h205: o_val = 'h7C12;
            'h206: o_val = 'h7B49;
            'h207: o_val = 'h7A80;
            'h208: o_val = 'h79B7;
            'h209: o_val = 'h78EE;
            'h20A: o_val = 'h7826;
            'h20B: o_val = 'h775D;
            'h20C: o_val = 'h7694;
            'h20D: o_val = 'h75CC;
            'h20E: o_val = 'h7504;
            'h20F: o_val = 'h743B;
            'h210: o_val = 'h7373;
            'h211: o_val = 'h72AB;
            'h212: o_val = 'h71E3;
            'h213: o_val = 'h711C;
            'h214: o_val = 'h7054;
            'h215: o_val = 'h6F8C;
            'h216: o_val = 'h6EC5;
            'h217: o_val = 'h6DFE;
            'h218: o_val = 'h6D37;
            'h219: o_val = 'h6C70;
            'h21A: o_val = 'h6BAA;
            'h21B: o_val = 'h6AE3;
            'h21C: o_val = 'h6A1D;
            'h21D: o_val = 'h6957;
            'h21E: o_val = 'h6891;
            'h21F: o_val = 'h67CC;
            'h220: o_val = 'h6706;
            'h221: o_val = 'h6641;
            'h222: o_val = 'h657C;
            'h223: o_val = 'h64B8;
            'h224: o_val = 'h63F4;
            'h225: o_val = 'h6330;
            'h226: o_val = 'h626C;
            'h227: o_val = 'h61A8;
            'h228: o_val = 'h60E5;
            'h229: o_val = 'h6022;
            'h22A: o_val = 'h5F60;
            'h22B: o_val = 'h5E9D;
            'h22C: o_val = 'h5DDB;
            'h22D: o_val = 'h5D1A;
            'h22E: o_val = 'h5C59;
            'h22F: o_val = 'h5B98;
            'h230: o_val = 'h5AD7;
            'h231: o_val = 'h5A17;
            'h232: o_val = 'h5957;
            'h233: o_val = 'h5898;
            'h234: o_val = 'h57D8;
            'h235: o_val = 'h571A;
            'h236: o_val = 'h565B;
            'h237: o_val = 'h559D;
            'h238: o_val = 'h54E0;
            'h239: o_val = 'h5423;
            'h23A: o_val = 'h5366;
            'h23B: o_val = 'h52AA;
            'h23C: o_val = 'h51EE;
            'h23D: o_val = 'h5133;
            'h23E: o_val = 'h5078;
            'h23F: o_val = 'h4FBD;
            'h240: o_val = 'h4F03;
            'h241: o_val = 'h4E4A;
            'h242: o_val = 'h4D91;
            'h243: o_val = 'h4CD8;
            'h244: o_val = 'h4C20;
            'h245: o_val = 'h4B69;
            'h246: o_val = 'h4AB2;
            'h247: o_val = 'h49FB;
            'h248: o_val = 'h4945;
            'h249: o_val = 'h4890;
            'h24A: o_val = 'h47DB;
            'h24B: o_val = 'h4726;
            'h24C: o_val = 'h4672;
            'h24D: o_val = 'h45BF;
            'h24E: o_val = 'h450C;
            'h24F: o_val = 'h445A;
            'h250: o_val = 'h43A9;
            'h251: o_val = 'h42F7;
            'h252: o_val = 'h4247;
            'h253: o_val = 'h4197;
            'h254: o_val = 'h40E8;
            'h255: o_val = 'h4039;
            'h256: o_val = 'h3F8B;
            'h257: o_val = 'h3EDE;
            'h258: o_val = 'h3E31;
            'h259: o_val = 'h3D85;
            'h25A: o_val = 'h3CDA;
            'h25B: o_val = 'h3C2F;
            'h25C: o_val = 'h3B84;
            'h25D: o_val = 'h3ADB;
            'h25E: o_val = 'h3A32;
            'h25F: o_val = 'h398A;
            'h260: o_val = 'h38E2;
            'h261: o_val = 'h383C;
            'h262: o_val = 'h3795;
            'h263: o_val = 'h36F0;
            'h264: o_val = 'h364B;
            'h265: o_val = 'h35A7;
            'h266: o_val = 'h3504;
            'h267: o_val = 'h3461;
            'h268: o_val = 'h33BF;
            'h269: o_val = 'h331E;
            'h26A: o_val = 'h327E;
            'h26B: o_val = 'h31DE;
            'h26C: o_val = 'h313F;
            'h26D: o_val = 'h30A1;
            'h26E: o_val = 'h3004;
            'h26F: o_val = 'h2F67;
            'h270: o_val = 'h2ECC;
            'h271: o_val = 'h2E30;
            'h272: o_val = 'h2D96;
            'h273: o_val = 'h2CFD;
            'h274: o_val = 'h2C64;
            'h275: o_val = 'h2BCC;
            'h276: o_val = 'h2B35;
            'h277: o_val = 'h2A9F;
            'h278: o_val = 'h2A0A;
            'h279: o_val = 'h2975;
            'h27A: o_val = 'h28E1;
            'h27B: o_val = 'h284F;
            'h27C: o_val = 'h27BC;
            'h27D: o_val = 'h272B;
            'h27E: o_val = 'h269B;
            'h27F: o_val = 'h260B;
            'h280: o_val = 'h257D;
            'h281: o_val = 'h24EF;
            'h282: o_val = 'h2462;
            'h283: o_val = 'h23D6;
            'h284: o_val = 'h234B;
            'h285: o_val = 'h22C1;
            'h286: o_val = 'h2238;
            'h287: o_val = 'h21AF;
            'h288: o_val = 'h2128;
            'h289: o_val = 'h20A1;
            'h28A: o_val = 'h201C;
            'h28B: o_val = 'h1F97;
            'h28C: o_val = 'h1F13;
            'h28D: o_val = 'h1E90;
            'h28E: o_val = 'h1E0E;
            'h28F: o_val = 'h1D8D;
            'h290: o_val = 'h1D0D;
            'h291: o_val = 'h1C8E;
            'h292: o_val = 'h1C10;
            'h293: o_val = 'h1B93;
            'h294: o_val = 'h1B17;
            'h295: o_val = 'h1A9C;
            'h296: o_val = 'h1A21;
            'h297: o_val = 'h19A8;
            'h298: o_val = 'h1930;
            'h299: o_val = 'h18B9;
            'h29A: o_val = 'h1842;
            'h29B: o_val = 'h17CD;
            'h29C: o_val = 'h1759;
            'h29D: o_val = 'h16E6;
            'h29E: o_val = 'h1673;
            'h29F: o_val = 'h1602;
            'h2A0: o_val = 'h1592;
            'h2A1: o_val = 'h1523;
            'h2A2: o_val = 'h14B4;
            'h2A3: o_val = 'h1447;
            'h2A4: o_val = 'h13DB;
            'h2A5: o_val = 'h1370;
            'h2A6: o_val = 'h1306;
            'h2A7: o_val = 'h129D;
            'h2A8: o_val = 'h1235;
            'h2A9: o_val = 'h11CF;
            'h2AA: o_val = 'h1169;
            'h2AB: o_val = 'h1104;
            'h2AC: o_val = 'h10A0;
            'h2AD: o_val = 'h103E;
            'h2AE: o_val = 'h0FDC;
            'h2AF: o_val = 'h0F7C;
            'h2B0: o_val = 'h0F1D;
            'h2B1: o_val = 'h0EBE;
            'h2B2: o_val = 'h0E61;
            'h2B3: o_val = 'h0E05;
            'h2B4: o_val = 'h0DAA;
            'h2B5: o_val = 'h0D50;
            'h2B6: o_val = 'h0CF8;
            'h2B7: o_val = 'h0CA0;
            'h2B8: o_val = 'h0C4A;
            'h2B9: o_val = 'h0BF4;
            'h2BA: o_val = 'h0BA0;
            'h2BB: o_val = 'h0B4D;
            'h2BC: o_val = 'h0AFB;
            'h2BD: o_val = 'h0AAA;
            'h2BE: o_val = 'h0A5A;
            'h2BF: o_val = 'h0A0B;
            'h2C0: o_val = 'h09BE;
            'h2C1: o_val = 'h0971;
            'h2C2: o_val = 'h0926;
            'h2C3: o_val = 'h08DC;
            'h2C4: o_val = 'h0893;
            'h2C5: o_val = 'h084B;
            'h2C6: o_val = 'h0805;
            'h2C7: o_val = 'h07BF;
            'h2C8: o_val = 'h077B;
            'h2C9: o_val = 'h0738;
            'h2CA: o_val = 'h06F6;
            'h2CB: o_val = 'h06B5;
            'h2CC: o_val = 'h0675;
            'h2CD: o_val = 'h0637;
            'h2CE: o_val = 'h05FA;
            'h2CF: o_val = 'h05BD;
            'h2D0: o_val = 'h0582;
            'h2D1: o_val = 'h0549;
            'h2D2: o_val = 'h0510;
            'h2D3: o_val = 'h04D9;
            'h2D4: o_val = 'h04A2;
            'h2D5: o_val = 'h046D;
            'h2D6: o_val = 'h043A;
            'h2D7: o_val = 'h0407;
            'h2D8: o_val = 'h03D6;
            'h2D9: o_val = 'h03A5;
            'h2DA: o_val = 'h0376;
            'h2DB: o_val = 'h0348;
            'h2DC: o_val = 'h031C;
            'h2DD: o_val = 'h02F0;
            'h2DE: o_val = 'h02C6;
            'h2DF: o_val = 'h029D;
            'h2E0: o_val = 'h0275;
            'h2E1: o_val = 'h024E;
            'h2E2: o_val = 'h0229;
            'h2E3: o_val = 'h0205;
            'h2E4: o_val = 'h01E2;
            'h2E5: o_val = 'h01C0;
            'h2E6: o_val = 'h01A0;
            'h2E7: o_val = 'h0180;
            'h2E8: o_val = 'h0162;
            'h2E9: o_val = 'h0145;
            'h2EA: o_val = 'h012A;
            'h2EB: o_val = 'h010F;
            'h2EC: o_val = 'h00F6;
            'h2ED: o_val = 'h00DE;
            'h2EE: o_val = 'h00C7;
            'h2EF: o_val = 'h00B2;
            'h2F0: o_val = 'h009D;
            'h2F1: o_val = 'h008A;
            'h2F2: o_val = 'h0078;
            'h2F3: o_val = 'h0068;
            'h2F4: o_val = 'h0058;
            'h2F5: o_val = 'h004A;
            'h2F6: o_val = 'h003D;
            'h2F7: o_val = 'h0031;
            'h2F8: o_val = 'h0027;
            'h2F9: o_val = 'h001E;
            'h2FA: o_val = 'h0016;
            'h2FB: o_val = 'h000F;
            'h2FC: o_val = 'h0009;
            'h2FD: o_val = 'h0005;
            'h2FE: o_val = 'h0002;
            'h2FF: o_val = 'h0000;
            'h300: o_val = 'h0000;
            'h301: o_val = 'h0000;
            'h302: o_val = 'h0002;
            'h303: o_val = 'h0005;
            'h304: o_val = 'h0009;
            'h305: o_val = 'h000F;
            'h306: o_val = 'h0016;
            'h307: o_val = 'h001E;
            'h308: o_val = 'h0027;
            'h309: o_val = 'h0031;
            'h30A: o_val = 'h003D;
            'h30B: o_val = 'h004A;
            'h30C: o_val = 'h0058;
            'h30D: o_val = 'h0068;
            'h30E: o_val = 'h0078;
            'h30F: o_val = 'h008A;
            'h310: o_val = 'h009D;
            'h311: o_val = 'h00B2;
            'h312: o_val = 'h00C7;
            'h313: o_val = 'h00DE;
            'h314: o_val = 'h00F6;
            'h315: o_val = 'h010F;
            'h316: o_val = 'h012A;
            'h317: o_val = 'h0145;
            'h318: o_val = 'h0162;
            'h319: o_val = 'h0180;
            'h31A: o_val = 'h01A0;
            'h31B: o_val = 'h01C0;
            'h31C: o_val = 'h01E2;
            'h31D: o_val = 'h0205;
            'h31E: o_val = 'h0229;
            'h31F: o_val = 'h024E;
            'h320: o_val = 'h0275;
            'h321: o_val = 'h029D;
            'h322: o_val = 'h02C6;
            'h323: o_val = 'h02F0;
            'h324: o_val = 'h031C;
            'h325: o_val = 'h0348;
            'h326: o_val = 'h0376;
            'h327: o_val = 'h03A5;
            'h328: o_val = 'h03D6;
            'h329: o_val = 'h0407;
            'h32A: o_val = 'h043A;
            'h32B: o_val = 'h046D;
            'h32C: o_val = 'h04A2;
            'h32D: o_val = 'h04D9;
            'h32E: o_val = 'h0510;
            'h32F: o_val = 'h0549;
            'h330: o_val = 'h0582;
            'h331: o_val = 'h05BD;
            'h332: o_val = 'h05FA;
            'h333: o_val = 'h0637;
            'h334: o_val = 'h0675;
            'h335: o_val = 'h06B5;
            'h336: o_val = 'h06F6;
            'h337: o_val = 'h0738;
            'h338: o_val = 'h077B;
            'h339: o_val = 'h07BF;
            'h33A: o_val = 'h0805;
            'h33B: o_val = 'h084B;
            'h33C: o_val = 'h0893;
            'h33D: o_val = 'h08DC;
            'h33E: o_val = 'h0926;
            'h33F: o_val = 'h0971;
            'h340: o_val = 'h09BE;
            'h341: o_val = 'h0A0B;
            'h342: o_val = 'h0A5A;
            'h343: o_val = 'h0AAA;
            'h344: o_val = 'h0AFB;
            'h345: o_val = 'h0B4D;
            'h346: o_val = 'h0BA0;
            'h347: o_val = 'h0BF4;
            'h348: o_val = 'h0C4A;
            'h349: o_val = 'h0CA0;
            'h34A: o_val = 'h0CF8;
            'h34B: o_val = 'h0D50;
            'h34C: o_val = 'h0DAA;
            'h34D: o_val = 'h0E05;
            'h34E: o_val = 'h0E61;
            'h34F: o_val = 'h0EBE;
            'h350: o_val = 'h0F1D;
            'h351: o_val = 'h0F7C;
            'h352: o_val = 'h0FDC;
            'h353: o_val = 'h103E;
            'h354: o_val = 'h10A0;
            'h355: o_val = 'h1104;
            'h356: o_val = 'h1169;
            'h357: o_val = 'h11CF;
            'h358: o_val = 'h1235;
            'h359: o_val = 'h129D;
            'h35A: o_val = 'h1306;
            'h35B: o_val = 'h1370;
            'h35C: o_val = 'h13DB;
            'h35D: o_val = 'h1447;
            'h35E: o_val = 'h14B4;
            'h35F: o_val = 'h1523;
            'h360: o_val = 'h1592;
            'h361: o_val = 'h1602;
            'h362: o_val = 'h1673;
            'h363: o_val = 'h16E6;
            'h364: o_val = 'h1759;
            'h365: o_val = 'h17CD;
            'h366: o_val = 'h1842;
            'h367: o_val = 'h18B9;
            'h368: o_val = 'h1930;
            'h369: o_val = 'h19A8;
            'h36A: o_val = 'h1A21;
            'h36B: o_val = 'h1A9C;
            'h36C: o_val = 'h1B17;
            'h36D: o_val = 'h1B93;
            'h36E: o_val = 'h1C10;
            'h36F: o_val = 'h1C8E;
            'h370: o_val = 'h1D0D;
            'h371: o_val = 'h1D8D;
            'h372: o_val = 'h1E0E;
            'h373: o_val = 'h1E90;
            'h374: o_val = 'h1F13;
            'h375: o_val = 'h1F97;
            'h376: o_val = 'h201C;
            'h377: o_val = 'h20A1;
            'h378: o_val = 'h2128;
            'h379: o_val = 'h21AF;
            'h37A: o_val = 'h2238;
            'h37B: o_val = 'h22C1;
            'h37C: o_val = 'h234B;
            'h37D: o_val = 'h23D6;
            'h37E: o_val = 'h2462;
            'h37F: o_val = 'h24EF;
            'h380: o_val = 'h257D;
            'h381: o_val = 'h260B;
            'h382: o_val = 'h269B;
            'h383: o_val = 'h272B;
            'h384: o_val = 'h27BC;
            'h385: o_val = 'h284F;
            'h386: o_val = 'h28E1;
            'h387: o_val = 'h2975;
            'h388: o_val = 'h2A0A;
            'h389: o_val = 'h2A9F;
            'h38A: o_val = 'h2B35;
            'h38B: o_val = 'h2BCC;
            'h38C: o_val = 'h2C64;
            'h38D: o_val = 'h2CFD;
            'h38E: o_val = 'h2D96;
            'h38F: o_val = 'h2E30;
            'h390: o_val = 'h2ECC;
            'h391: o_val = 'h2F67;
            'h392: o_val = 'h3004;
            'h393: o_val = 'h30A1;
            'h394: o_val = 'h313F;
            'h395: o_val = 'h31DE;
            'h396: o_val = 'h327E;
            'h397: o_val = 'h331E;
            'h398: o_val = 'h33BF;
            'h399: o_val = 'h3461;
            'h39A: o_val = 'h3504;
            'h39B: o_val = 'h35A7;
            'h39C: o_val = 'h364B;
            'h39D: o_val = 'h36F0;
            'h39E: o_val = 'h3795;
            'h39F: o_val = 'h383C;
            'h3A0: o_val = 'h38E2;
            'h3A1: o_val = 'h398A;
            'h3A2: o_val = 'h3A32;
            'h3A3: o_val = 'h3ADB;
            'h3A4: o_val = 'h3B84;
            'h3A5: o_val = 'h3C2F;
            'h3A6: o_val = 'h3CDA;
            'h3A7: o_val = 'h3D85;
            'h3A8: o_val = 'h3E31;
            'h3A9: o_val = 'h3EDE;
            'h3AA: o_val = 'h3F8B;
            'h3AB: o_val = 'h4039;
            'h3AC: o_val = 'h40E8;
            'h3AD: o_val = 'h4197;
            'h3AE: o_val = 'h4247;
            'h3AF: o_val = 'h42F7;
            'h3B0: o_val = 'h43A9;
            'h3B1: o_val = 'h445A;
            'h3B2: o_val = 'h450C;
            'h3B3: o_val = 'h45BF;
            'h3B4: o_val = 'h4672;
            'h3B5: o_val = 'h4726;
            'h3B6: o_val = 'h47DB;
            'h3B7: o_val = 'h4890;
            'h3B8: o_val = 'h4945;
            'h3B9: o_val = 'h49FB;
            'h3BA: o_val = 'h4AB2;
            'h3BB: o_val = 'h4B69;
            'h3BC: o_val = 'h4C20;
            'h3BD: o_val = 'h4CD8;
            'h3BE: o_val = 'h4D91;
            'h3BF: o_val = 'h4E4A;
            'h3C0: o_val = 'h4F03;
            'h3C1: o_val = 'h4FBD;
            'h3C2: o_val = 'h5078;
            'h3C3: o_val = 'h5133;
            'h3C4: o_val = 'h51EE;
            'h3C5: o_val = 'h52AA;
            'h3C6: o_val = 'h5366;
            'h3C7: o_val = 'h5423;
            'h3C8: o_val = 'h54E0;
            'h3C9: o_val = 'h559D;
            'h3CA: o_val = 'h565B;
            'h3CB: o_val = 'h571A;
            'h3CC: o_val = 'h57D8;
            'h3CD: o_val = 'h5898;
            'h3CE: o_val = 'h5957;
            'h3CF: o_val = 'h5A17;
            'h3D0: o_val = 'h5AD7;
            'h3D1: o_val = 'h5B98;
            'h3D2: o_val = 'h5C59;
            'h3D3: o_val = 'h5D1A;
            'h3D4: o_val = 'h5DDB;
            'h3D5: o_val = 'h5E9D;
            'h3D6: o_val = 'h5F60;
            'h3D7: o_val = 'h6022;
            'h3D8: o_val = 'h60E5;
            'h3D9: o_val = 'h61A8;
            'h3DA: o_val = 'h626C;
            'h3DB: o_val = 'h6330;
            'h3DC: o_val = 'h63F4;
            'h3DD: o_val = 'h64B8;
            'h3DE: o_val = 'h657C;
            'h3DF: o_val = 'h6641;
            'h3E0: o_val = 'h6706;
            'h3E1: o_val = 'h67CC;
            'h3E2: o_val = 'h6891;
            'h3E3: o_val = 'h6957;
            'h3E4: o_val = 'h6A1D;
            'h3E5: o_val = 'h6AE3;
            'h3E6: o_val = 'h6BAA;
            'h3E7: o_val = 'h6C70;
            'h3E8: o_val = 'h6D37;
            'h3E9: o_val = 'h6DFE;
            'h3EA: o_val = 'h6EC5;
            'h3EB: o_val = 'h6F8C;
            'h3EC: o_val = 'h7054;
            'h3ED: o_val = 'h711C;
            'h3EE: o_val = 'h71E3;
            'h3EF: o_val = 'h72AB;
            'h3F0: o_val = 'h7373;
            'h3F1: o_val = 'h743B;
            'h3F2: o_val = 'h7504;
            'h3F3: o_val = 'h75CC;
            'h3F4: o_val = 'h7694;
            'h3F5: o_val = 'h775D;
            'h3F6: o_val = 'h7826;
            'h3F7: o_val = 'h78EE;
            'h3F8: o_val = 'h79B7;
            'h3F9: o_val = 'h7A80;
            'h3FA: o_val = 'h7B49;
            'h3FB: o_val = 'h7C12;
            'h3FC: o_val = 'h7CDB;
            'h3FD: o_val = 'h7DA4;
            'h3FE: o_val = 'h7E6D;
            'h3FF: o_val = 'h7F36;
        endcase
    end
endmodule