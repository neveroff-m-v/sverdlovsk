/*
    SVERDLOVSK
    system verilog library

    Neveroff M.V.
    2025
*/

/// Статистика по тестированию (тестбенчу)
package testbench;

/// Тип ошибки
class error_type;
endclass

/// Отчет о испытании
class report;
endclass

/// Отчет о тестировании (тестбенче)
class testbench;
endclass

endpackage 
