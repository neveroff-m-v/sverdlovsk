package const;

class const;

    static const int pulldown = 0;
    static const int pullup = 1;

endclass

endpackage