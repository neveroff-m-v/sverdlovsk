package constant;

class pull;

    static int down = 0;
    static int up = 1;

endclass

endpackage