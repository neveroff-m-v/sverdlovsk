// Таблица COS (10'b -> 16'b)
module ram_cos (
    i_val,
    o_val
    );

    input  [15:0] i_val;
    output [15:0] o_val;

    always_comb begin
        o_val = 'h0000;

        case (i_val[15:6])
            'h000: o_val = 'hFFFF;
            'h001: o_val = 'hFFFE;
            'h002: o_val = 'hFFFC;
            'h003: o_val = 'hFFF9;
            'h004: o_val = 'hFFF5;
            'h005: o_val = 'hFFEF;
            'h006: o_val = 'hFFE8;
            'h007: o_val = 'hFFE0;
            'h008: o_val = 'hFFD7;
            'h009: o_val = 'hFFCD;
            'h00A: o_val = 'hFFC1;
            'h00B: o_val = 'hFFB4;
            'h00C: o_val = 'hFFA6;
            'h00D: o_val = 'hFF96;
            'h00E: o_val = 'hFF86;
            'h00F: o_val = 'hFF74;
            'h010: o_val = 'hFF61;
            'h011: o_val = 'hFF4C;
            'h012: o_val = 'hFF37;
            'h013: o_val = 'hFF20;
            'h014: o_val = 'hFF08;
            'h015: o_val = 'hFEEF;
            'h016: o_val = 'hFED4;
            'h017: o_val = 'hFEB9;
            'h018: o_val = 'hFE9C;
            'h019: o_val = 'hFE7E;
            'h01A: o_val = 'hFE5E;
            'h01B: o_val = 'hFE3E;
            'h01C: o_val = 'hFE1C;
            'h01D: o_val = 'hFDF9;
            'h01E: o_val = 'hFDD5;
            'h01F: o_val = 'hFDB0;
            'h020: o_val = 'hFD89;
            'h021: o_val = 'hFD61;
            'h022: o_val = 'hFD38;
            'h023: o_val = 'hFD0E;
            'h024: o_val = 'hFCE2;
            'h025: o_val = 'hFCB6;
            'h026: o_val = 'hFC88;
            'h027: o_val = 'hFC59;
            'h028: o_val = 'hFC28;
            'h029: o_val = 'hFBF7;
            'h02A: o_val = 'hFBC4;
            'h02B: o_val = 'hFB91;
            'h02C: o_val = 'hFB5C;
            'h02D: o_val = 'hFB25;
            'h02E: o_val = 'hFAEE;
            'h02F: o_val = 'hFAB5;
            'h030: o_val = 'hFA7C;
            'h031: o_val = 'hFA41;
            'h032: o_val = 'hFA04;
            'h033: o_val = 'hF9C7;
            'h034: o_val = 'hF989;
            'h035: o_val = 'hF949;
            'h036: o_val = 'hF908;
            'h037: o_val = 'hF8C6;
            'h038: o_val = 'hF883;
            'h039: o_val = 'hF83F;
            'h03A: o_val = 'hF7F9;
            'h03B: o_val = 'hF7B3;
            'h03C: o_val = 'hF76B;
            'h03D: o_val = 'hF722;
            'h03E: o_val = 'hF6D8;
            'h03F: o_val = 'hF68D;
            'h040: o_val = 'hF640;
            'h041: o_val = 'hF5F3;
            'h042: o_val = 'hF5A4;
            'h043: o_val = 'hF554;
            'h044: o_val = 'hF503;
            'h045: o_val = 'hF4B1;
            'h046: o_val = 'hF45E;
            'h047: o_val = 'hF40A;
            'h048: o_val = 'hF3B4;
            'h049: o_val = 'hF35E;
            'h04A: o_val = 'hF306;
            'h04B: o_val = 'hF2AE;
            'h04C: o_val = 'hF254;
            'h04D: o_val = 'hF1F9;
            'h04E: o_val = 'hF19D;
            'h04F: o_val = 'hF140;
            'h050: o_val = 'hF0E1;
            'h051: o_val = 'hF082;
            'h052: o_val = 'hF022;
            'h053: o_val = 'hEFC0;
            'h054: o_val = 'hEF5E;
            'h055: o_val = 'hEEFA;
            'h056: o_val = 'hEE95;
            'h057: o_val = 'hEE2F;
            'h058: o_val = 'hEDC9;
            'h059: o_val = 'hED61;
            'h05A: o_val = 'hECF8;
            'h05B: o_val = 'hEC8E;
            'h05C: o_val = 'hEC23;
            'h05D: o_val = 'hEBB7;
            'h05E: o_val = 'hEB4A;
            'h05F: o_val = 'hEADB;
            'h060: o_val = 'hEA6C;
            'h061: o_val = 'hE9FC;
            'h062: o_val = 'hE98B;
            'h063: o_val = 'hE918;
            'h064: o_val = 'hE8A5;
            'h065: o_val = 'hE831;
            'h066: o_val = 'hE7BC;
            'h067: o_val = 'hE745;
            'h068: o_val = 'hE6CE;
            'h069: o_val = 'hE656;
            'h06A: o_val = 'hE5DD;
            'h06B: o_val = 'hE562;
            'h06C: o_val = 'hE4E7;
            'h06D: o_val = 'hE46B;
            'h06E: o_val = 'hE3EE;
            'h06F: o_val = 'hE370;
            'h070: o_val = 'hE2F1;
            'h071: o_val = 'hE271;
            'h072: o_val = 'hE1F0;
            'h073: o_val = 'hE16E;
            'h074: o_val = 'hE0EB;
            'h075: o_val = 'hE067;
            'h076: o_val = 'hDFE2;
            'h077: o_val = 'hDF5D;
            'h078: o_val = 'hDED6;
            'h079: o_val = 'hDE4F;
            'h07A: o_val = 'hDDC6;
            'h07B: o_val = 'hDD3D;
            'h07C: o_val = 'hDCB3;
            'h07D: o_val = 'hDC28;
            'h07E: o_val = 'hDB9C;
            'h07F: o_val = 'hDB0F;
            'h080: o_val = 'hDA81;
            'h081: o_val = 'hD9F3;
            'h082: o_val = 'hD963;
            'h083: o_val = 'hD8D3;
            'h084: o_val = 'hD842;
            'h085: o_val = 'hD7AF;
            'h086: o_val = 'hD71D;
            'h087: o_val = 'hD689;
            'h088: o_val = 'hD5F4;
            'h089: o_val = 'hD55F;
            'h08A: o_val = 'hD4C9;
            'h08B: o_val = 'hD432;
            'h08C: o_val = 'hD39A;
            'h08D: o_val = 'hD301;
            'h08E: o_val = 'hD268;
            'h08F: o_val = 'hD1CE;
            'h090: o_val = 'hD132;
            'h091: o_val = 'hD097;
            'h092: o_val = 'hCFFA;
            'h093: o_val = 'hCF5D;
            'h094: o_val = 'hCEBF;
            'h095: o_val = 'hCE20;
            'h096: o_val = 'hCD80;
            'h097: o_val = 'hCCE0;
            'h098: o_val = 'hCC3F;
            'h099: o_val = 'hCB9D;
            'h09A: o_val = 'hCAFA;
            'h09B: o_val = 'hCA57;
            'h09C: o_val = 'hC9B3;
            'h09D: o_val = 'hC90E;
            'h09E: o_val = 'hC869;
            'h09F: o_val = 'hC7C2;
            'h0A0: o_val = 'hC71C;
            'h0A1: o_val = 'hC674;
            'h0A2: o_val = 'hC5CC;
            'h0A3: o_val = 'hC523;
            'h0A4: o_val = 'hC47A;
            'h0A5: o_val = 'hC3CF;
            'h0A6: o_val = 'hC324;
            'h0A7: o_val = 'hC279;
            'h0A8: o_val = 'hC1CD;
            'h0A9: o_val = 'hC120;
            'h0AA: o_val = 'hC073;
            'h0AB: o_val = 'hBFC5;
            'h0AC: o_val = 'hBF16;
            'h0AD: o_val = 'hBE67;
            'h0AE: o_val = 'hBDB7;
            'h0AF: o_val = 'hBD07;
            'h0B0: o_val = 'hBC55;
            'h0B1: o_val = 'hBBA4;
            'h0B2: o_val = 'hBAF2;
            'h0B3: o_val = 'hBA3F;
            'h0B4: o_val = 'hB98C;
            'h0B5: o_val = 'hB8D8;
            'h0B6: o_val = 'hB823;
            'h0B7: o_val = 'hB76E;
            'h0B8: o_val = 'hB6B9;
            'h0B9: o_val = 'hB603;
            'h0BA: o_val = 'hB54C;
            'h0BB: o_val = 'hB495;
            'h0BC: o_val = 'hB3DE;
            'h0BD: o_val = 'hB326;
            'h0BE: o_val = 'hB26D;
            'h0BF: o_val = 'hB1B4;
            'h0C0: o_val = 'hB0FB;
            'h0C1: o_val = 'hB041;
            'h0C2: o_val = 'hAF86;
            'h0C3: o_val = 'hAECB;
            'h0C4: o_val = 'hAE10;
            'h0C5: o_val = 'hAD54;
            'h0C6: o_val = 'hAC98;
            'h0C7: o_val = 'hABDB;
            'h0C8: o_val = 'hAB1E;
            'h0C9: o_val = 'hAA61;
            'h0CA: o_val = 'hA9A3;
            'h0CB: o_val = 'hA8E4;
            'h0CC: o_val = 'hA826;
            'h0CD: o_val = 'hA766;
            'h0CE: o_val = 'hA6A7;
            'h0CF: o_val = 'hA5E7;
            'h0D0: o_val = 'hA527;
            'h0D1: o_val = 'hA466;
            'h0D2: o_val = 'hA3A5;
            'h0D3: o_val = 'hA2E4;
            'h0D4: o_val = 'hA223;
            'h0D5: o_val = 'hA161;
            'h0D6: o_val = 'hA09E;
            'h0D7: o_val = 'h9FDC;
            'h0D8: o_val = 'h9F19;
            'h0D9: o_val = 'h9E56;
            'h0DA: o_val = 'h9D92;
            'h0DB: o_val = 'h9CCE;
            'h0DC: o_val = 'h9C0A;
            'h0DD: o_val = 'h9B46;
            'h0DE: o_val = 'h9A82;
            'h0DF: o_val = 'h99BD;
            'h0E0: o_val = 'h98F8;
            'h0E1: o_val = 'h9832;
            'h0E2: o_val = 'h976D;
            'h0E3: o_val = 'h96A7;
            'h0E4: o_val = 'h95E1;
            'h0E5: o_val = 'h951B;
            'h0E6: o_val = 'h9454;
            'h0E7: o_val = 'h938E;
            'h0E8: o_val = 'h92C7;
            'h0E9: o_val = 'h9200;
            'h0EA: o_val = 'h9139;
            'h0EB: o_val = 'h9072;
            'h0EC: o_val = 'h8FAA;
            'h0ED: o_val = 'h8EE2;
            'h0EE: o_val = 'h8E1B;
            'h0EF: o_val = 'h8D53;
            'h0F0: o_val = 'h8C8B;
            'h0F1: o_val = 'h8BC3;
            'h0F2: o_val = 'h8AFA;
            'h0F3: o_val = 'h8A32;
            'h0F4: o_val = 'h896A;
            'h0F5: o_val = 'h88A1;
            'h0F6: o_val = 'h87D8;
            'h0F7: o_val = 'h8710;
            'h0F8: o_val = 'h8647;
            'h0F9: o_val = 'h857E;
            'h0FA: o_val = 'h84B5;
            'h0FB: o_val = 'h83EC;
            'h0FC: o_val = 'h8323;
            'h0FD: o_val = 'h825A;
            'h0FE: o_val = 'h8191;
            'h0FF: o_val = 'h80C8;
            'h100: o_val = 'h7FFF;
            'h101: o_val = 'h7F36;
            'h102: o_val = 'h7E6D;
            'h103: o_val = 'h7DA4;
            'h104: o_val = 'h7CDB;
            'h105: o_val = 'h7C12;
            'h106: o_val = 'h7B49;
            'h107: o_val = 'h7A80;
            'h108: o_val = 'h79B7;
            'h109: o_val = 'h78EE;
            'h10A: o_val = 'h7826;
            'h10B: o_val = 'h775D;
            'h10C: o_val = 'h7694;
            'h10D: o_val = 'h75CC;
            'h10E: o_val = 'h7504;
            'h10F: o_val = 'h743B;
            'h110: o_val = 'h7373;
            'h111: o_val = 'h72AB;
            'h112: o_val = 'h71E3;
            'h113: o_val = 'h711C;
            'h114: o_val = 'h7054;
            'h115: o_val = 'h6F8C;
            'h116: o_val = 'h6EC5;
            'h117: o_val = 'h6DFE;
            'h118: o_val = 'h6D37;
            'h119: o_val = 'h6C70;
            'h11A: o_val = 'h6BAA;
            'h11B: o_val = 'h6AE3;
            'h11C: o_val = 'h6A1D;
            'h11D: o_val = 'h6957;
            'h11E: o_val = 'h6891;
            'h11F: o_val = 'h67CC;
            'h120: o_val = 'h6706;
            'h121: o_val = 'h6641;
            'h122: o_val = 'h657C;
            'h123: o_val = 'h64B8;
            'h124: o_val = 'h63F4;
            'h125: o_val = 'h6330;
            'h126: o_val = 'h626C;
            'h127: o_val = 'h61A8;
            'h128: o_val = 'h60E5;
            'h129: o_val = 'h6022;
            'h12A: o_val = 'h5F60;
            'h12B: o_val = 'h5E9D;
            'h12C: o_val = 'h5DDB;
            'h12D: o_val = 'h5D1A;
            'h12E: o_val = 'h5C59;
            'h12F: o_val = 'h5B98;
            'h130: o_val = 'h5AD7;
            'h131: o_val = 'h5A17;
            'h132: o_val = 'h5957;
            'h133: o_val = 'h5898;
            'h134: o_val = 'h57D8;
            'h135: o_val = 'h571A;
            'h136: o_val = 'h565B;
            'h137: o_val = 'h559D;
            'h138: o_val = 'h54E0;
            'h139: o_val = 'h5423;
            'h13A: o_val = 'h5366;
            'h13B: o_val = 'h52AA;
            'h13C: o_val = 'h51EE;
            'h13D: o_val = 'h5133;
            'h13E: o_val = 'h5078;
            'h13F: o_val = 'h4FBD;
            'h140: o_val = 'h4F03;
            'h141: o_val = 'h4E4A;
            'h142: o_val = 'h4D91;
            'h143: o_val = 'h4CD8;
            'h144: o_val = 'h4C20;
            'h145: o_val = 'h4B69;
            'h146: o_val = 'h4AB2;
            'h147: o_val = 'h49FB;
            'h148: o_val = 'h4945;
            'h149: o_val = 'h4890;
            'h14A: o_val = 'h47DB;
            'h14B: o_val = 'h4726;
            'h14C: o_val = 'h4672;
            'h14D: o_val = 'h45BF;
            'h14E: o_val = 'h450C;
            'h14F: o_val = 'h445A;
            'h150: o_val = 'h43A9;
            'h151: o_val = 'h42F7;
            'h152: o_val = 'h4247;
            'h153: o_val = 'h4197;
            'h154: o_val = 'h40E8;
            'h155: o_val = 'h4039;
            'h156: o_val = 'h3F8B;
            'h157: o_val = 'h3EDE;
            'h158: o_val = 'h3E31;
            'h159: o_val = 'h3D85;
            'h15A: o_val = 'h3CDA;
            'h15B: o_val = 'h3C2F;
            'h15C: o_val = 'h3B84;
            'h15D: o_val = 'h3ADB;
            'h15E: o_val = 'h3A32;
            'h15F: o_val = 'h398A;
            'h160: o_val = 'h38E2;
            'h161: o_val = 'h383C;
            'h162: o_val = 'h3795;
            'h163: o_val = 'h36F0;
            'h164: o_val = 'h364B;
            'h165: o_val = 'h35A7;
            'h166: o_val = 'h3504;
            'h167: o_val = 'h3461;
            'h168: o_val = 'h33BF;
            'h169: o_val = 'h331E;
            'h16A: o_val = 'h327E;
            'h16B: o_val = 'h31DE;
            'h16C: o_val = 'h313F;
            'h16D: o_val = 'h30A1;
            'h16E: o_val = 'h3004;
            'h16F: o_val = 'h2F67;
            'h170: o_val = 'h2ECC;
            'h171: o_val = 'h2E30;
            'h172: o_val = 'h2D96;
            'h173: o_val = 'h2CFD;
            'h174: o_val = 'h2C64;
            'h175: o_val = 'h2BCC;
            'h176: o_val = 'h2B35;
            'h177: o_val = 'h2A9F;
            'h178: o_val = 'h2A0A;
            'h179: o_val = 'h2975;
            'h17A: o_val = 'h28E1;
            'h17B: o_val = 'h284F;
            'h17C: o_val = 'h27BC;
            'h17D: o_val = 'h272B;
            'h17E: o_val = 'h269B;
            'h17F: o_val = 'h260B;
            'h180: o_val = 'h257D;
            'h181: o_val = 'h24EF;
            'h182: o_val = 'h2462;
            'h183: o_val = 'h23D6;
            'h184: o_val = 'h234B;
            'h185: o_val = 'h22C1;
            'h186: o_val = 'h2238;
            'h187: o_val = 'h21AF;
            'h188: o_val = 'h2128;
            'h189: o_val = 'h20A1;
            'h18A: o_val = 'h201C;
            'h18B: o_val = 'h1F97;
            'h18C: o_val = 'h1F13;
            'h18D: o_val = 'h1E90;
            'h18E: o_val = 'h1E0E;
            'h18F: o_val = 'h1D8D;
            'h190: o_val = 'h1D0D;
            'h191: o_val = 'h1C8E;
            'h192: o_val = 'h1C10;
            'h193: o_val = 'h1B93;
            'h194: o_val = 'h1B17;
            'h195: o_val = 'h1A9C;
            'h196: o_val = 'h1A21;
            'h197: o_val = 'h19A8;
            'h198: o_val = 'h1930;
            'h199: o_val = 'h18B9;
            'h19A: o_val = 'h1842;
            'h19B: o_val = 'h17CD;
            'h19C: o_val = 'h1759;
            'h19D: o_val = 'h16E6;
            'h19E: o_val = 'h1673;
            'h19F: o_val = 'h1602;
            'h1A0: o_val = 'h1592;
            'h1A1: o_val = 'h1523;
            'h1A2: o_val = 'h14B4;
            'h1A3: o_val = 'h1447;
            'h1A4: o_val = 'h13DB;
            'h1A5: o_val = 'h1370;
            'h1A6: o_val = 'h1306;
            'h1A7: o_val = 'h129D;
            'h1A8: o_val = 'h1235;
            'h1A9: o_val = 'h11CF;
            'h1AA: o_val = 'h1169;
            'h1AB: o_val = 'h1104;
            'h1AC: o_val = 'h10A0;
            'h1AD: o_val = 'h103E;
            'h1AE: o_val = 'h0FDC;
            'h1AF: o_val = 'h0F7C;
            'h1B0: o_val = 'h0F1D;
            'h1B1: o_val = 'h0EBE;
            'h1B2: o_val = 'h0E61;
            'h1B3: o_val = 'h0E05;
            'h1B4: o_val = 'h0DAA;
            'h1B5: o_val = 'h0D50;
            'h1B6: o_val = 'h0CF8;
            'h1B7: o_val = 'h0CA0;
            'h1B8: o_val = 'h0C4A;
            'h1B9: o_val = 'h0BF4;
            'h1BA: o_val = 'h0BA0;
            'h1BB: o_val = 'h0B4D;
            'h1BC: o_val = 'h0AFB;
            'h1BD: o_val = 'h0AAA;
            'h1BE: o_val = 'h0A5A;
            'h1BF: o_val = 'h0A0B;
            'h1C0: o_val = 'h09BE;
            'h1C1: o_val = 'h0971;
            'h1C2: o_val = 'h0926;
            'h1C3: o_val = 'h08DC;
            'h1C4: o_val = 'h0893;
            'h1C5: o_val = 'h084B;
            'h1C6: o_val = 'h0805;
            'h1C7: o_val = 'h07BF;
            'h1C8: o_val = 'h077B;
            'h1C9: o_val = 'h0738;
            'h1CA: o_val = 'h06F6;
            'h1CB: o_val = 'h06B5;
            'h1CC: o_val = 'h0675;
            'h1CD: o_val = 'h0637;
            'h1CE: o_val = 'h05FA;
            'h1CF: o_val = 'h05BD;
            'h1D0: o_val = 'h0582;
            'h1D1: o_val = 'h0549;
            'h1D2: o_val = 'h0510;
            'h1D3: o_val = 'h04D9;
            'h1D4: o_val = 'h04A2;
            'h1D5: o_val = 'h046D;
            'h1D6: o_val = 'h043A;
            'h1D7: o_val = 'h0407;
            'h1D8: o_val = 'h03D6;
            'h1D9: o_val = 'h03A5;
            'h1DA: o_val = 'h0376;
            'h1DB: o_val = 'h0348;
            'h1DC: o_val = 'h031C;
            'h1DD: o_val = 'h02F0;
            'h1DE: o_val = 'h02C6;
            'h1DF: o_val = 'h029D;
            'h1E0: o_val = 'h0275;
            'h1E1: o_val = 'h024E;
            'h1E2: o_val = 'h0229;
            'h1E3: o_val = 'h0205;
            'h1E4: o_val = 'h01E2;
            'h1E5: o_val = 'h01C0;
            'h1E6: o_val = 'h01A0;
            'h1E7: o_val = 'h0180;
            'h1E8: o_val = 'h0162;
            'h1E9: o_val = 'h0145;
            'h1EA: o_val = 'h012A;
            'h1EB: o_val = 'h010F;
            'h1EC: o_val = 'h00F6;
            'h1ED: o_val = 'h00DE;
            'h1EE: o_val = 'h00C7;
            'h1EF: o_val = 'h00B2;
            'h1F0: o_val = 'h009D;
            'h1F1: o_val = 'h008A;
            'h1F2: o_val = 'h0078;
            'h1F3: o_val = 'h0068;
            'h1F4: o_val = 'h0058;
            'h1F5: o_val = 'h004A;
            'h1F6: o_val = 'h003D;
            'h1F7: o_val = 'h0031;
            'h1F8: o_val = 'h0027;
            'h1F9: o_val = 'h001E;
            'h1FA: o_val = 'h0016;
            'h1FB: o_val = 'h000F;
            'h1FC: o_val = 'h0009;
            'h1FD: o_val = 'h0005;
            'h1FE: o_val = 'h0002;
            'h1FF: o_val = 'h0000;
            'h200: o_val = 'h0000;
            'h201: o_val = 'h0000;
            'h202: o_val = 'h0002;
            'h203: o_val = 'h0005;
            'h204: o_val = 'h0009;
            'h205: o_val = 'h000F;
            'h206: o_val = 'h0016;
            'h207: o_val = 'h001E;
            'h208: o_val = 'h0027;
            'h209: o_val = 'h0031;
            'h20A: o_val = 'h003D;
            'h20B: o_val = 'h004A;
            'h20C: o_val = 'h0058;
            'h20D: o_val = 'h0068;
            'h20E: o_val = 'h0078;
            'h20F: o_val = 'h008A;
            'h210: o_val = 'h009D;
            'h211: o_val = 'h00B2;
            'h212: o_val = 'h00C7;
            'h213: o_val = 'h00DE;
            'h214: o_val = 'h00F6;
            'h215: o_val = 'h010F;
            'h216: o_val = 'h012A;
            'h217: o_val = 'h0145;
            'h218: o_val = 'h0162;
            'h219: o_val = 'h0180;
            'h21A: o_val = 'h01A0;
            'h21B: o_val = 'h01C0;
            'h21C: o_val = 'h01E2;
            'h21D: o_val = 'h0205;
            'h21E: o_val = 'h0229;
            'h21F: o_val = 'h024E;
            'h220: o_val = 'h0275;
            'h221: o_val = 'h029D;
            'h222: o_val = 'h02C6;
            'h223: o_val = 'h02F0;
            'h224: o_val = 'h031C;
            'h225: o_val = 'h0348;
            'h226: o_val = 'h0376;
            'h227: o_val = 'h03A5;
            'h228: o_val = 'h03D6;
            'h229: o_val = 'h0407;
            'h22A: o_val = 'h043A;
            'h22B: o_val = 'h046D;
            'h22C: o_val = 'h04A2;
            'h22D: o_val = 'h04D9;
            'h22E: o_val = 'h0510;
            'h22F: o_val = 'h0549;
            'h230: o_val = 'h0582;
            'h231: o_val = 'h05BD;
            'h232: o_val = 'h05FA;
            'h233: o_val = 'h0637;
            'h234: o_val = 'h0675;
            'h235: o_val = 'h06B5;
            'h236: o_val = 'h06F6;
            'h237: o_val = 'h0738;
            'h238: o_val = 'h077B;
            'h239: o_val = 'h07BF;
            'h23A: o_val = 'h0805;
            'h23B: o_val = 'h084B;
            'h23C: o_val = 'h0893;
            'h23D: o_val = 'h08DC;
            'h23E: o_val = 'h0926;
            'h23F: o_val = 'h0971;
            'h240: o_val = 'h09BE;
            'h241: o_val = 'h0A0B;
            'h242: o_val = 'h0A5A;
            'h243: o_val = 'h0AAA;
            'h244: o_val = 'h0AFB;
            'h245: o_val = 'h0B4D;
            'h246: o_val = 'h0BA0;
            'h247: o_val = 'h0BF4;
            'h248: o_val = 'h0C4A;
            'h249: o_val = 'h0CA0;
            'h24A: o_val = 'h0CF8;
            'h24B: o_val = 'h0D50;
            'h24C: o_val = 'h0DAA;
            'h24D: o_val = 'h0E05;
            'h24E: o_val = 'h0E61;
            'h24F: o_val = 'h0EBE;
            'h250: o_val = 'h0F1D;
            'h251: o_val = 'h0F7C;
            'h252: o_val = 'h0FDC;
            'h253: o_val = 'h103E;
            'h254: o_val = 'h10A0;
            'h255: o_val = 'h1104;
            'h256: o_val = 'h1169;
            'h257: o_val = 'h11CF;
            'h258: o_val = 'h1235;
            'h259: o_val = 'h129D;
            'h25A: o_val = 'h1306;
            'h25B: o_val = 'h1370;
            'h25C: o_val = 'h13DB;
            'h25D: o_val = 'h1447;
            'h25E: o_val = 'h14B4;
            'h25F: o_val = 'h1523;
            'h260: o_val = 'h1592;
            'h261: o_val = 'h1602;
            'h262: o_val = 'h1673;
            'h263: o_val = 'h16E6;
            'h264: o_val = 'h1759;
            'h265: o_val = 'h17CD;
            'h266: o_val = 'h1842;
            'h267: o_val = 'h18B9;
            'h268: o_val = 'h1930;
            'h269: o_val = 'h19A8;
            'h26A: o_val = 'h1A21;
            'h26B: o_val = 'h1A9C;
            'h26C: o_val = 'h1B17;
            'h26D: o_val = 'h1B93;
            'h26E: o_val = 'h1C10;
            'h26F: o_val = 'h1C8E;
            'h270: o_val = 'h1D0D;
            'h271: o_val = 'h1D8D;
            'h272: o_val = 'h1E0E;
            'h273: o_val = 'h1E90;
            'h274: o_val = 'h1F13;
            'h275: o_val = 'h1F97;
            'h276: o_val = 'h201C;
            'h277: o_val = 'h20A1;
            'h278: o_val = 'h2128;
            'h279: o_val = 'h21AF;
            'h27A: o_val = 'h2238;
            'h27B: o_val = 'h22C1;
            'h27C: o_val = 'h234B;
            'h27D: o_val = 'h23D6;
            'h27E: o_val = 'h2462;
            'h27F: o_val = 'h24EF;
            'h280: o_val = 'h257D;
            'h281: o_val = 'h260B;
            'h282: o_val = 'h269B;
            'h283: o_val = 'h272B;
            'h284: o_val = 'h27BC;
            'h285: o_val = 'h284F;
            'h286: o_val = 'h28E1;
            'h287: o_val = 'h2975;
            'h288: o_val = 'h2A0A;
            'h289: o_val = 'h2A9F;
            'h28A: o_val = 'h2B35;
            'h28B: o_val = 'h2BCC;
            'h28C: o_val = 'h2C64;
            'h28D: o_val = 'h2CFD;
            'h28E: o_val = 'h2D96;
            'h28F: o_val = 'h2E30;
            'h290: o_val = 'h2ECC;
            'h291: o_val = 'h2F67;
            'h292: o_val = 'h3004;
            'h293: o_val = 'h30A1;
            'h294: o_val = 'h313F;
            'h295: o_val = 'h31DE;
            'h296: o_val = 'h327E;
            'h297: o_val = 'h331E;
            'h298: o_val = 'h33BF;
            'h299: o_val = 'h3461;
            'h29A: o_val = 'h3504;
            'h29B: o_val = 'h35A7;
            'h29C: o_val = 'h364B;
            'h29D: o_val = 'h36F0;
            'h29E: o_val = 'h3795;
            'h29F: o_val = 'h383C;
            'h2A0: o_val = 'h38E2;
            'h2A1: o_val = 'h398A;
            'h2A2: o_val = 'h3A32;
            'h2A3: o_val = 'h3ADB;
            'h2A4: o_val = 'h3B84;
            'h2A5: o_val = 'h3C2F;
            'h2A6: o_val = 'h3CDA;
            'h2A7: o_val = 'h3D85;
            'h2A8: o_val = 'h3E31;
            'h2A9: o_val = 'h3EDE;
            'h2AA: o_val = 'h3F8B;
            'h2AB: o_val = 'h4039;
            'h2AC: o_val = 'h40E8;
            'h2AD: o_val = 'h4197;
            'h2AE: o_val = 'h4247;
            'h2AF: o_val = 'h42F7;
            'h2B0: o_val = 'h43A9;
            'h2B1: o_val = 'h445A;
            'h2B2: o_val = 'h450C;
            'h2B3: o_val = 'h45BF;
            'h2B4: o_val = 'h4672;
            'h2B5: o_val = 'h4726;
            'h2B6: o_val = 'h47DB;
            'h2B7: o_val = 'h4890;
            'h2B8: o_val = 'h4945;
            'h2B9: o_val = 'h49FB;
            'h2BA: o_val = 'h4AB2;
            'h2BB: o_val = 'h4B69;
            'h2BC: o_val = 'h4C20;
            'h2BD: o_val = 'h4CD8;
            'h2BE: o_val = 'h4D91;
            'h2BF: o_val = 'h4E4A;
            'h2C0: o_val = 'h4F03;
            'h2C1: o_val = 'h4FBD;
            'h2C2: o_val = 'h5078;
            'h2C3: o_val = 'h5133;
            'h2C4: o_val = 'h51EE;
            'h2C5: o_val = 'h52AA;
            'h2C6: o_val = 'h5366;
            'h2C7: o_val = 'h5423;
            'h2C8: o_val = 'h54E0;
            'h2C9: o_val = 'h559D;
            'h2CA: o_val = 'h565B;
            'h2CB: o_val = 'h571A;
            'h2CC: o_val = 'h57D8;
            'h2CD: o_val = 'h5898;
            'h2CE: o_val = 'h5957;
            'h2CF: o_val = 'h5A17;
            'h2D0: o_val = 'h5AD7;
            'h2D1: o_val = 'h5B98;
            'h2D2: o_val = 'h5C59;
            'h2D3: o_val = 'h5D1A;
            'h2D4: o_val = 'h5DDB;
            'h2D5: o_val = 'h5E9D;
            'h2D6: o_val = 'h5F60;
            'h2D7: o_val = 'h6022;
            'h2D8: o_val = 'h60E5;
            'h2D9: o_val = 'h61A8;
            'h2DA: o_val = 'h626C;
            'h2DB: o_val = 'h6330;
            'h2DC: o_val = 'h63F4;
            'h2DD: o_val = 'h64B8;
            'h2DE: o_val = 'h657C;
            'h2DF: o_val = 'h6641;
            'h2E0: o_val = 'h6706;
            'h2E1: o_val = 'h67CC;
            'h2E2: o_val = 'h6891;
            'h2E3: o_val = 'h6957;
            'h2E4: o_val = 'h6A1D;
            'h2E5: o_val = 'h6AE3;
            'h2E6: o_val = 'h6BAA;
            'h2E7: o_val = 'h6C70;
            'h2E8: o_val = 'h6D37;
            'h2E9: o_val = 'h6DFE;
            'h2EA: o_val = 'h6EC5;
            'h2EB: o_val = 'h6F8C;
            'h2EC: o_val = 'h7054;
            'h2ED: o_val = 'h711C;
            'h2EE: o_val = 'h71E3;
            'h2EF: o_val = 'h72AB;
            'h2F0: o_val = 'h7373;
            'h2F1: o_val = 'h743B;
            'h2F2: o_val = 'h7504;
            'h2F3: o_val = 'h75CC;
            'h2F4: o_val = 'h7694;
            'h2F5: o_val = 'h775D;
            'h2F6: o_val = 'h7826;
            'h2F7: o_val = 'h78EE;
            'h2F8: o_val = 'h79B7;
            'h2F9: o_val = 'h7A80;
            'h2FA: o_val = 'h7B49;
            'h2FB: o_val = 'h7C12;
            'h2FC: o_val = 'h7CDB;
            'h2FD: o_val = 'h7DA4;
            'h2FE: o_val = 'h7E6D;
            'h2FF: o_val = 'h7F36;
            'h300: o_val = 'h7FFF;
            'h301: o_val = 'h80C8;
            'h302: o_val = 'h8191;
            'h303: o_val = 'h825A;
            'h304: o_val = 'h8323;
            'h305: o_val = 'h83EC;
            'h306: o_val = 'h84B5;
            'h307: o_val = 'h857E;
            'h308: o_val = 'h8647;
            'h309: o_val = 'h8710;
            'h30A: o_val = 'h87D8;
            'h30B: o_val = 'h88A1;
            'h30C: o_val = 'h896A;
            'h30D: o_val = 'h8A32;
            'h30E: o_val = 'h8AFA;
            'h30F: o_val = 'h8BC3;
            'h310: o_val = 'h8C8B;
            'h311: o_val = 'h8D53;
            'h312: o_val = 'h8E1B;
            'h313: o_val = 'h8EE2;
            'h314: o_val = 'h8FAA;
            'h315: o_val = 'h9072;
            'h316: o_val = 'h9139;
            'h317: o_val = 'h9200;
            'h318: o_val = 'h92C7;
            'h319: o_val = 'h938E;
            'h31A: o_val = 'h9454;
            'h31B: o_val = 'h951B;
            'h31C: o_val = 'h95E1;
            'h31D: o_val = 'h96A7;
            'h31E: o_val = 'h976D;
            'h31F: o_val = 'h9832;
            'h320: o_val = 'h98F8;
            'h321: o_val = 'h99BD;
            'h322: o_val = 'h9A82;
            'h323: o_val = 'h9B46;
            'h324: o_val = 'h9C0A;
            'h325: o_val = 'h9CCE;
            'h326: o_val = 'h9D92;
            'h327: o_val = 'h9E56;
            'h328: o_val = 'h9F19;
            'h329: o_val = 'h9FDC;
            'h32A: o_val = 'hA09E;
            'h32B: o_val = 'hA161;
            'h32C: o_val = 'hA223;
            'h32D: o_val = 'hA2E4;
            'h32E: o_val = 'hA3A5;
            'h32F: o_val = 'hA466;
            'h330: o_val = 'hA527;
            'h331: o_val = 'hA5E7;
            'h332: o_val = 'hA6A7;
            'h333: o_val = 'hA766;
            'h334: o_val = 'hA826;
            'h335: o_val = 'hA8E4;
            'h336: o_val = 'hA9A3;
            'h337: o_val = 'hAA61;
            'h338: o_val = 'hAB1E;
            'h339: o_val = 'hABDB;
            'h33A: o_val = 'hAC98;
            'h33B: o_val = 'hAD54;
            'h33C: o_val = 'hAE10;
            'h33D: o_val = 'hAECB;
            'h33E: o_val = 'hAF86;
            'h33F: o_val = 'hB041;
            'h340: o_val = 'hB0FB;
            'h341: o_val = 'hB1B4;
            'h342: o_val = 'hB26D;
            'h343: o_val = 'hB326;
            'h344: o_val = 'hB3DE;
            'h345: o_val = 'hB495;
            'h346: o_val = 'hB54C;
            'h347: o_val = 'hB603;
            'h348: o_val = 'hB6B9;
            'h349: o_val = 'hB76E;
            'h34A: o_val = 'hB823;
            'h34B: o_val = 'hB8D8;
            'h34C: o_val = 'hB98C;
            'h34D: o_val = 'hBA3F;
            'h34E: o_val = 'hBAF2;
            'h34F: o_val = 'hBBA4;
            'h350: o_val = 'hBC55;
            'h351: o_val = 'hBD07;
            'h352: o_val = 'hBDB7;
            'h353: o_val = 'hBE67;
            'h354: o_val = 'hBF16;
            'h355: o_val = 'hBFC5;
            'h356: o_val = 'hC073;
            'h357: o_val = 'hC120;
            'h358: o_val = 'hC1CD;
            'h359: o_val = 'hC279;
            'h35A: o_val = 'hC324;
            'h35B: o_val = 'hC3CF;
            'h35C: o_val = 'hC47A;
            'h35D: o_val = 'hC523;
            'h35E: o_val = 'hC5CC;
            'h35F: o_val = 'hC674;
            'h360: o_val = 'hC71C;
            'h361: o_val = 'hC7C2;
            'h362: o_val = 'hC869;
            'h363: o_val = 'hC90E;
            'h364: o_val = 'hC9B3;
            'h365: o_val = 'hCA57;
            'h366: o_val = 'hCAFA;
            'h367: o_val = 'hCB9D;
            'h368: o_val = 'hCC3F;
            'h369: o_val = 'hCCE0;
            'h36A: o_val = 'hCD80;
            'h36B: o_val = 'hCE20;
            'h36C: o_val = 'hCEBF;
            'h36D: o_val = 'hCF5D;
            'h36E: o_val = 'hCFFA;
            'h36F: o_val = 'hD097;
            'h370: o_val = 'hD132;
            'h371: o_val = 'hD1CE;
            'h372: o_val = 'hD268;
            'h373: o_val = 'hD301;
            'h374: o_val = 'hD39A;
            'h375: o_val = 'hD432;
            'h376: o_val = 'hD4C9;
            'h377: o_val = 'hD55F;
            'h378: o_val = 'hD5F4;
            'h379: o_val = 'hD689;
            'h37A: o_val = 'hD71D;
            'h37B: o_val = 'hD7AF;
            'h37C: o_val = 'hD842;
            'h37D: o_val = 'hD8D3;
            'h37E: o_val = 'hD963;
            'h37F: o_val = 'hD9F3;
            'h380: o_val = 'hDA81;
            'h381: o_val = 'hDB0F;
            'h382: o_val = 'hDB9C;
            'h383: o_val = 'hDC28;
            'h384: o_val = 'hDCB3;
            'h385: o_val = 'hDD3D;
            'h386: o_val = 'hDDC6;
            'h387: o_val = 'hDE4F;
            'h388: o_val = 'hDED6;
            'h389: o_val = 'hDF5D;
            'h38A: o_val = 'hDFE2;
            'h38B: o_val = 'hE067;
            'h38C: o_val = 'hE0EB;
            'h38D: o_val = 'hE16E;
            'h38E: o_val = 'hE1F0;
            'h38F: o_val = 'hE271;
            'h390: o_val = 'hE2F1;
            'h391: o_val = 'hE370;
            'h392: o_val = 'hE3EE;
            'h393: o_val = 'hE46B;
            'h394: o_val = 'hE4E7;
            'h395: o_val = 'hE562;
            'h396: o_val = 'hE5DD;
            'h397: o_val = 'hE656;
            'h398: o_val = 'hE6CE;
            'h399: o_val = 'hE745;
            'h39A: o_val = 'hE7BC;
            'h39B: o_val = 'hE831;
            'h39C: o_val = 'hE8A5;
            'h39D: o_val = 'hE918;
            'h39E: o_val = 'hE98B;
            'h39F: o_val = 'hE9FC;
            'h3A0: o_val = 'hEA6C;
            'h3A1: o_val = 'hEADB;
            'h3A2: o_val = 'hEB4A;
            'h3A3: o_val = 'hEBB7;
            'h3A4: o_val = 'hEC23;
            'h3A5: o_val = 'hEC8E;
            'h3A6: o_val = 'hECF8;
            'h3A7: o_val = 'hED61;
            'h3A8: o_val = 'hEDC9;
            'h3A9: o_val = 'hEE2F;
            'h3AA: o_val = 'hEE95;
            'h3AB: o_val = 'hEEFA;
            'h3AC: o_val = 'hEF5E;
            'h3AD: o_val = 'hEFC0;
            'h3AE: o_val = 'hF022;
            'h3AF: o_val = 'hF082;
            'h3B0: o_val = 'hF0E1;
            'h3B1: o_val = 'hF140;
            'h3B2: o_val = 'hF19D;
            'h3B3: o_val = 'hF1F9;
            'h3B4: o_val = 'hF254;
            'h3B5: o_val = 'hF2AE;
            'h3B6: o_val = 'hF306;
            'h3B7: o_val = 'hF35E;
            'h3B8: o_val = 'hF3B4;
            'h3B9: o_val = 'hF40A;
            'h3BA: o_val = 'hF45E;
            'h3BB: o_val = 'hF4B1;
            'h3BC: o_val = 'hF503;
            'h3BD: o_val = 'hF554;
            'h3BE: o_val = 'hF5A4;
            'h3BF: o_val = 'hF5F3;
            'h3C0: o_val = 'hF640;
            'h3C1: o_val = 'hF68D;
            'h3C2: o_val = 'hF6D8;
            'h3C3: o_val = 'hF722;
            'h3C4: o_val = 'hF76B;
            'h3C5: o_val = 'hF7B3;
            'h3C6: o_val = 'hF7F9;
            'h3C7: o_val = 'hF83F;
            'h3C8: o_val = 'hF883;
            'h3C9: o_val = 'hF8C6;
            'h3CA: o_val = 'hF908;
            'h3CB: o_val = 'hF949;
            'h3CC: o_val = 'hF989;
            'h3CD: o_val = 'hF9C7;
            'h3CE: o_val = 'hFA04;
            'h3CF: o_val = 'hFA41;
            'h3D0: o_val = 'hFA7C;
            'h3D1: o_val = 'hFAB5;
            'h3D2: o_val = 'hFAEE;
            'h3D3: o_val = 'hFB25;
            'h3D4: o_val = 'hFB5C;
            'h3D5: o_val = 'hFB91;
            'h3D6: o_val = 'hFBC4;
            'h3D7: o_val = 'hFBF7;
            'h3D8: o_val = 'hFC28;
            'h3D9: o_val = 'hFC59;
            'h3DA: o_val = 'hFC88;
            'h3DB: o_val = 'hFCB6;
            'h3DC: o_val = 'hFCE2;
            'h3DD: o_val = 'hFD0E;
            'h3DE: o_val = 'hFD38;
            'h3DF: o_val = 'hFD61;
            'h3E0: o_val = 'hFD89;
            'h3E1: o_val = 'hFDB0;
            'h3E2: o_val = 'hFDD5;
            'h3E3: o_val = 'hFDF9;
            'h3E4: o_val = 'hFE1C;
            'h3E5: o_val = 'hFE3E;
            'h3E6: o_val = 'hFE5E;
            'h3E7: o_val = 'hFE7E;
            'h3E8: o_val = 'hFE9C;
            'h3E9: o_val = 'hFEB9;
            'h3EA: o_val = 'hFED4;
            'h3EB: o_val = 'hFEEF;
            'h3EC: o_val = 'hFF08;
            'h3ED: o_val = 'hFF20;
            'h3EE: o_val = 'hFF37;
            'h3EF: o_val = 'hFF4C;
            'h3F0: o_val = 'hFF61;
            'h3F1: o_val = 'hFF74;
            'h3F2: o_val = 'hFF86;
            'h3F3: o_val = 'hFF96;
            'h3F4: o_val = 'hFFA6;
            'h3F5: o_val = 'hFFB4;
            'h3F6: o_val = 'hFFC1;
            'h3F7: o_val = 'hFFCD;
            'h3F8: o_val = 'hFFD7;
            'h3F9: o_val = 'hFFE0;
            'h3FA: o_val = 'hFFE8;
            'h3FB: o_val = 'hFFEF;
            'h3FC: o_val = 'hFFF5;
            'h3FD: o_val = 'hFFF9;
            'h3FE: o_val = 'hFFFC;
            'h3FF: o_val = 'hFFFE;
        endcase
    end
endmodule